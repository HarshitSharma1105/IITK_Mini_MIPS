module FPU(input float,input[31:0] instruction,input cc);


always @(posedge float)

    $display("Float");



endmodule